.subckt PC817 1 2 3 4

* Node 1 -> DA
* Node 2 -> DK
* Node 3 -> QE
* Node 4 -> QC
* Node 5 -> QB

DIN 1 6 dmodel
VT 6 2 0
CIO 1 4 1e-12
QOUT 4 5 3 qmodel
RFX 3 5 1e9
BFX 3 5 I=0+0.00091067*I(VT)+1.2307*I(VT)*I(VT)
RB  5  3 1meg

* Default values used in dmodel:
*   TT=0 BV=infinite

.MODEL dmodel d
+IS=1.4174e-12 RS=1.77049 N=1.96012 XTI=4
+EG=1.50946 CJO=1e-11 VJ=0.75 M=0.5 FC=0.5
.MODEL qmodel npn
+IS=2.04341e-10 BF=1000 NF=1.04784 VAF=74.9441
+IKF=0.0207989 ISE=1e-08 NE=4 BR=0.1
+NR=1.5 VAR=1.1341 IKR=0.207989 ISC=9.99193e-14
+NC=2.00279 RB=10 IRB=0.2 RBM=10
+RE=4.57626 RC=100 XTB=0.1 XTI=2.77723 EG=0.1
+CJE=9.76772e-12 VJE=0.4 MJE=0.180481 TF=1.00004e-09
+XTF=1 VTF=10 ITF=0.01 CJC=1.96829e-11
+VJC=0.59397 MJC=0.415235 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1

.ends PC817

* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt MC33076  1 2 3 4 5
*
  c1   11 12 11.72E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 6.063E6 -1E3 1E3 6E6 -6E6
  ga    6  0 11 12 659.7E-6
  gcm   0  6 10 99 20.86E-9
  iee   3 10 dc 78.20E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   4 11 1.516E3
  rc2   4 12 1.516E3
  re1  13 10 850.4
  re2  14 10 850.4
  ree  10 99 2.558E6
  ro1   8  5 50
  ro2   7 99 50
  rp    3  4 10.89E3
  vb    9  0 dc 0
  vc    3 53 dc 1.200
  ve   54  4 dc 1.200
  vlim  7  8 dc 0
  vlp  91  0 dc 250
  vln   0 92 dc 250
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx PNP(Is=800.0E-18 Bf=390)
.ends

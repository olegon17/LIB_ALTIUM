********************************************************************
*
*  Copyright (c) International Rectifier
*
*  IR2113: High and Low Side Driver
*   
*  Ports 
*    VDD: Logic Supply
*    HIN: Logic Input for High Side Gate Driver Output(HO), in phase
*    SD:  Logic Input for Shutdown
*    LIN: Logic Input for Low Side Gate Driver Output(LO), in phase
*    VSS: Logic Ground
*    VB:  High Side Floating Supply 
*    HO:  High Side Gate Diver Output
*    VS:  High Side Floating Supply Return
*    VCC: Low Side Supply
*    LO:  Low Side Gate Driver Output
*    COM: Low Side Return
*
*  Created by Pspice Version 8 
*
*  Date Created: 03/25/2003
*
********************************************************************
*
*  This behavioral model was developed in compliance with Data Sheet 
*  No. PD60147-R except noted below: 
*  (1) There is no frequency effect on temperature.
*  (2) The power dissipation is different. 
*  (3) The values of output high/low short circuit current are adjusted 
*      for the proper modeling of turn-on rise/turn-off fall time.
*  (4) The "Low side return (COM)" pin must be grounded.
*
***********************************************************************

.SUBCKT IR2113 VDD HIN SD LIN VSS HO VB VS VCC COM LO 
+PARAMS:  
+         T1=-40 T2=25 T3=125
+         V1=10 V2=15 V3=20
+         tonT1=90n tonT2=120n tonT3=170n
+         tonV1=140n tonV2=120n tonV3=100n
+         toffT1=77n toffT2=94n toffT3=130n
+         toffV1=115n toffV2=94n toffV3=75n
+         tonVdd1=125n tonVdd2=120n tonVdd3=115n
+         toffVdd1=113n toffVdd2=94n toffVdd3=72n

.MODEL diode25 d
+IS=1.0e-14 RS=0.01 N=1 EG=1.11
+XTI=3 BV=25 IBV=0.0001 CJO=0
+VJ=0.75 M=0.333 FC=0.5 TT=0
+KF=0 AF=1

.MODEL diode625 d
+IS=1.0e-14 RS=0.01 N=1 EG=1.11
+XTI=3 BV=625 IBV=0.0001 CJO=0
+VJ=0.75 M=0.333 FC=0.5 TT=0
+KF=0 AF=1

C_MD1_C2         VSS MD2_Nor3b_2  10p  
C_MD1_C3         VSS MD2_Inv2_1  10p  
C_MD1_C1         VSS MD2_Inv1_1  1n  
D_MD1_D2         VSS HIN diode25 
D_MD1_D3         SD VDD diode25 
D_MD1_D4         VSS SD diode25 
D_MD1_D5         LIN VDD diode25 
D_MD1_D6         VSS LIN diode25 
D_MD1_D7         VSS VDD diode25 
D_MD1_D1         HIN VDD diode25 
C_MD1_Trig3_CTrig         VSS MD2_Inv2_1  10p  
R_MD1_Trig3_R1Trig         MD1_Trig3_3 VDD  100Meg  
R_MD1_Trig3_R2Trig         MD1_Trig3_4 MD1_Trig3_3  66.7Meg  
R_MD1_Trig3_R3Trig         VSS MD1_Trig3_4  106.1Meg  
X_MD1_Trig3_Comp         LIN MD1_Trig3_3 MD2_Inv2_1 com COMP
S_MD1_Trig3_PTrig         MD1_Trig3_4 VSS MD2_Inv2_1 VSS _MD1_Trig3_PTrig
RS_MD1_Trig3_PTrig        MD2_Inv2_1 VSS 1G
.MODEL        _MD1_Trig3_PTrig VSWITCH Roff=1e9 Ron=1 Voff=0.01 Von=4.99
R_MD1_R1         VSS HIN 750k TC=-0.00783811, 0.0000372046
R_MD1_R2         VSS SD 750k TC=-0.00783811, 0.0000372046
C_MD1_Trig1_CTrig         VSS MD2_Inv1_1  10p  
R_MD1_Trig1_R1Trig         MD1_Trig1_3 VDD  100Meg  
R_MD1_Trig1_R2Trig         MD1_Trig1_4 MD1_Trig1_3  66.7Meg  
R_MD1_Trig1_R3Trig         VSS MD1_Trig1_4  106.1Meg  
X_MD1_Trig1_Comp         HIN MD1_Trig1_3 MD2_Inv1_1 com COMP
S_MD1_Trig1_PTrig         MD1_Trig1_4 VSS MD2_Inv1_1 VSS _MD1_Trig1_PTrig
RS_MD1_Trig1_PTrig        MD2_Inv1_1 VSS 1G
.MODEL        _MD1_Trig1_PTrig VSWITCH Roff=1e9 Ron=1 Voff=0.01 Von=4.99
C_MD1_Trig2_CTrig         VSS MD2_Nor3b_2  10p  
R_MD1_Trig2_R1Trig         MD1_Trig2_3 VDD  100Meg  
R_MD1_Trig2_R2Trig         MD1_Trig2_4 MD1_Trig2_3  66.7Meg  
R_MD1_Trig2_R3Trig         VSS MD1_Trig2_4  106.1Meg  
X_MD1_Trig2_Comp         SD MD1_Trig2_3 MD2_Nor3b_2 com COMP
S_MD1_Trig2_PTrig         MD1_Trig2_4 VSS MD2_Nor3b_2 VSS _MD1_Trig2_PTrig
RS_MD1_Trig2_PTrig        MD2_Nor3b_2 VSS 1G
.MODEL        _MD1_Trig2_PTrig VSWITCH Roff=1e9 Ron=1 Voff=0.01 Von=4.99
R_MD1_R3         VSS LIN 750k TC=-0.00783811, 0.0000372046
R_MD1_R4         VSS VDD 7.5Meg TC=-0.00505291, 0.0000236999
C_MD2_C1         VSS MD3_DlyHS_2  10p IC=0 
C_MD2_C2         VSS MD3_DlyLS_2  10p IC=0 
V_MD2_Inv1_V         MD2_Inv1_2 VSS 5V
C_MD2_Inv1_C         VSS MD2_Nor3a_3  1p  
S_MD2_Inv1_P         MD2_Inv1_2 MD2_Nor3a_3 MD2_Inv1_1 VSS _MD2_Inv1_P
RS_MD2_Inv1_P        MD2_Inv1_1 VSS 1G
.MODEL        _MD2_Inv1_P VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD2_Inv1_N         MD2_Nor3a_3 VSS MD2_Inv1_1 VSS _MD2_Inv1_N
RS_MD2_Inv1_N        MD2_Inv1_1 VSS 1G
.MODEL        _MD2_Inv1_N VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
V_MD2_Inv2_V         MD2_Inv2_2 VSS 5V
C_MD2_Inv2_C         VSS MD2_Nor3b_1  1p  
S_MD2_Inv2_P         MD2_Inv2_2 MD2_Nor3b_1 MD2_Inv2_1 VSS _MD2_Inv2_P
RS_MD2_Inv2_P        MD2_Inv2_1 VSS 1G
.MODEL        _MD2_Inv2_P VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD2_Inv2_N         MD2_Nor3b_1 VSS MD2_Inv2_1 VSS _MD2_Inv2_N
RS_MD2_Inv2_N        MD2_Inv2_1 VSS 1G
.MODEL        _MD2_Inv2_N VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
C_MD2_RS1_C7         MD2_RS1_6 MD2_RS1_5  10p  
C_MD2_RS1_C2         VSS MD2_Nor3a_3  10p IC=0 
C_MD2_RS1_C3         VSS MD2_Nor3b_2  10p IC=0 
C_MD2_RS1_C10         MD2_RS1_7 MD2_RS1_5  10p  
C_MD2_RS1_C11         MD2_RS1_3 MD2_RS1_7  10p  
C_MD2_RS1_C12         VSS MD2_RS1_3  10p  
C_MD2_RS1_C9         VSS MD2_Nor3a_1  10p  
C_MD2_RS1_C8         MD2_Nor3a_1 MD2_RS1_6  10p  
C_MD2_RS1_C1         VSS MD2_Nor3a_1  10p IC=0 
S_MD2_RS1_P1         MD2_RS1_5 MD2_RS1_6 MD2_Nor3a_3 VSS _MD2_RS1_P1
RS_MD2_RS1_P1        MD2_Nor3a_3 VSS 1G
.MODEL        _MD2_RS1_P1 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD2_RS1_P2         MD2_RS1_6 MD2_Nor3a_1 MD2_RS1_3 VSS _MD2_RS1_P2
RS_MD2_RS1_P2        MD2_RS1_3 VSS 1G
.MODEL        _MD2_RS1_P2 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD2_RS1_N1         MD2_Nor3a_1 VSS MD2_RS1_3 VSS _MD2_RS1_N1
RS_MD2_RS1_N1        MD2_RS1_3 VSS 1G
.MODEL        _MD2_RS1_N1 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
S_MD2_RS1_P3         MD2_RS1_5 MD2_RS1_7 MD2_Nor3b_2 VSS _MD2_RS1_P3
RS_MD2_RS1_P3        MD2_Nor3b_2 VSS 1G
.MODEL        _MD2_RS1_P3 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD2_RS1_P4         MD2_RS1_7 MD2_RS1_3 MD2_Nor3a_1 VSS _MD2_RS1_P4
RS_MD2_RS1_P4        MD2_Nor3a_1 VSS 1G
.MODEL        _MD2_RS1_P4 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD2_RS1_N3         MD2_RS1_3 VSS MD2_Nor3b_2 VSS _MD2_RS1_N3
RS_MD2_RS1_N3        MD2_Nor3b_2 VSS 1G
.MODEL        _MD2_RS1_N3 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
V_MD2_RS1_V1         MD2_RS1_5 VSS 5V
S_MD2_RS1_N4         MD2_RS1_3 VSS MD2_Nor3a_1 VSS _MD2_RS1_N4
RS_MD2_RS1_N4        MD2_Nor3a_1 VSS 1G
.MODEL        _MD2_RS1_N4 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
S_MD2_RS1_N2         MD2_Nor3a_1 VSS MD2_Nor3a_3 VSS _MD2_RS1_N2
RS_MD2_RS1_N2        MD2_Nor3a_3 VSS 1G
.MODEL        _MD2_RS1_N2 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
C_MD2_RS2_C7         MD2_RS2_6 MD2_RS2_5  10p  
C_MD2_RS2_C2         VSS MD2_Nor3b_1  10p IC=0 
C_MD2_RS2_C3         VSS MD2_Nor3b_2  10p IC=0 
C_MD2_RS2_C10         MD2_RS2_7 MD2_RS2_5  10p  
C_MD2_RS2_C11         MD2_RS2_3 MD2_RS2_7  10p  
C_MD2_RS2_C12         VSS MD2_RS2_3  10p  
C_MD2_RS2_C9         VSS MD2_Nor3b_3  10p  
C_MD2_RS2_C8         MD2_Nor3b_3 MD2_RS2_6  10p  
C_MD2_RS2_C1         VSS MD2_Nor3b_3  10p IC=0 
S_MD2_RS2_P1         MD2_RS2_5 MD2_RS2_6 MD2_Nor3b_1 VSS _MD2_RS2_P1
RS_MD2_RS2_P1        MD2_Nor3b_1 VSS 1G
.MODEL        _MD2_RS2_P1 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD2_RS2_P2         MD2_RS2_6 MD2_Nor3b_3 MD2_RS2_3 VSS _MD2_RS2_P2
RS_MD2_RS2_P2        MD2_RS2_3 VSS 1G
.MODEL        _MD2_RS2_P2 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD2_RS2_N1         MD2_Nor3b_3 VSS MD2_RS2_3 VSS _MD2_RS2_N1
RS_MD2_RS2_N1        MD2_RS2_3 VSS 1G
.MODEL        _MD2_RS2_N1 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
S_MD2_RS2_P3         MD2_RS2_5 MD2_RS2_7 MD2_Nor3b_2 VSS _MD2_RS2_P3
RS_MD2_RS2_P3        MD2_Nor3b_2 VSS 1G
.MODEL        _MD2_RS2_P3 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD2_RS2_P4         MD2_RS2_7 MD2_RS2_3 MD2_Nor3b_3 VSS _MD2_RS2_P4
RS_MD2_RS2_P4        MD2_Nor3b_3 VSS 1G
.MODEL        _MD2_RS2_P4 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD2_RS2_N3         MD2_RS2_3 VSS MD2_Nor3b_2 VSS _MD2_RS2_N3
RS_MD2_RS2_N3        MD2_Nor3b_2 VSS 1G
.MODEL        _MD2_RS2_N3 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
V_MD2_RS2_V1         MD2_RS2_5 VSS 5V
S_MD2_RS2_N4         MD2_RS2_3 VSS MD2_Nor3b_3 VSS _MD2_RS2_N4
RS_MD2_RS2_N4        MD2_Nor3b_3 VSS 1G
.MODEL        _MD2_RS2_N4 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
S_MD2_RS2_N2         MD2_Nor3b_3 VSS MD2_Nor3b_1 VSS _MD2_RS2_N2
RS_MD2_RS2_N2        MD2_Nor3b_1 VSS 1G
.MODEL        _MD2_RS2_N2 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
S_MD2_Nor3a_P1         MD2_Nor3a_4 MD2_Nor3a_5 MD2_Nor3a_1 VSS _MD2_Nor3a_P1
RS_MD2_Nor3a_P1        MD2_Nor3a_1 VSS 1G
.MODEL        _MD2_Nor3a_P1 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD2_Nor3a_P2         MD2_Nor3a_5 MD2_Nor3a_6 MD2_Nor3b_2 VSS _MD2_Nor3a_P2
RS_MD2_Nor3a_P2        MD2_Nor3b_2 VSS 1G
.MODEL        _MD2_Nor3a_P2 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD2_Nor3a_P3         MD2_Nor3a_6 MD3_DlyHS_2 MD2_Nor3a_3 VSS _MD2_Nor3a_P3
RS_MD2_Nor3a_P3        MD2_Nor3a_3 VSS 1G
.MODEL        _MD2_Nor3a_P3 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD2_Nor3a_N1         MD3_DlyHS_2 VSS MD2_Nor3b_2 VSS _MD2_Nor3a_N1
RS_MD2_Nor3a_N1        MD2_Nor3b_2 VSS 1G
.MODEL        _MD2_Nor3a_N1 VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
V_MD2_Nor3a_V         MD2_Nor3a_4 VSS 5V
S_MD2_Nor3a_N2         MD3_DlyHS_2 VSS MD2_Nor3a_1 VSS _MD2_Nor3a_N2
RS_MD2_Nor3a_N2        MD2_Nor3a_1 VSS 1G
.MODEL        _MD2_Nor3a_N2 VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
S_MD2_Nor3a_N3         MD3_DlyHS_2 VSS MD2_Nor3a_3 VSS _MD2_Nor3a_N3
RS_MD2_Nor3a_N3        MD2_Nor3a_3 VSS 1G
.MODEL        _MD2_Nor3a_N3 VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
S_MD2_Nor3b_P1         MD2_Nor3b_4 MD2_Nor3b_5 MD2_Nor3b_1 VSS _MD2_Nor3b_P1
RS_MD2_Nor3b_P1        MD2_Nor3b_1 VSS 1G
.MODEL        _MD2_Nor3b_P1 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD2_Nor3b_P2         MD2_Nor3b_5 MD2_Nor3b_6 MD2_Nor3b_2 VSS _MD2_Nor3b_P2
RS_MD2_Nor3b_P2        MD2_Nor3b_2 VSS 1G
.MODEL        _MD2_Nor3b_P2 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD2_Nor3b_P3         MD2_Nor3b_6 MD3_DlyLS_2 MD2_Nor3b_3 VSS _MD2_Nor3b_P3
RS_MD2_Nor3b_P3        MD2_Nor3b_3 VSS 1G
.MODEL        _MD2_Nor3b_P3 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD2_Nor3b_N1         MD3_DlyLS_2 VSS MD2_Nor3b_2 VSS _MD2_Nor3b_N1
RS_MD2_Nor3b_N1        MD2_Nor3b_2 VSS 1G
.MODEL        _MD2_Nor3b_N1 VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
V_MD2_Nor3b_V         MD2_Nor3b_4 VSS 5V
S_MD2_Nor3b_N2         MD3_DlyLS_2 VSS MD2_Nor3b_1 VSS _MD2_Nor3b_N2
RS_MD2_Nor3b_N2        MD2_Nor3b_1 VSS 1G
.MODEL        _MD2_Nor3b_N2 VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
S_MD2_Nor3b_N3         MD3_DlyLS_2 VSS MD2_Nor3b_3 VSS _MD2_Nor3b_N3
RS_MD2_Nor3b_N3        MD2_Nor3b_3 VSS 1G
.MODEL        _MD2_Nor3b_N3 VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
D_MD5_D2         com LO diode25 
D_MD5_D1         LO VCC diode25 
C_MD5_C         com LO  10p  
C_MD5_Uvcc_c1         MD5_Uvcc_2 MD5_Uvcc_3  10n  
C_MD5_Uvcc_c2         MD5_Uvcc_4 MD5_Uvcc_2  10n  
C_MD5_Uvcc_c3         com MD4_Inv5_1  10p  
E_MD5_Uvcc_ABM2         MD5_Uvcc_3 com   VALUE { 8.3+(8.8-8.3)/(125+40)*(TEMP+40)  
+   }
E_MD5_Uvcc_ABM3         MD5_Uvcc_4 com   VALUE { 8.0+(8.5-8.0)/(125+40)*(TEMP+40)  
+   }
X_MD5_Uvcc_Comp         VCC MD5_Uvcc_2 MD4_Inv5_1 com COMP
S_MD5_Uvcc_P         MD5_Uvcc_3 MD5_Uvcc_2 MD4_Inv5_1 com _MD5_Uvcc_P
RS_MD5_Uvcc_P        MD4_Inv5_1 com 1G
.MODEL        _MD5_Uvcc_P VSWITCH Roff=1e6 Ron=1 Voff=4.99 Von=0.01
S_MD5_Uvcc_N         MD5_Uvcc_2 MD5_Uvcc_4 MD4_Inv5_1 com _MD5_Uvcc_N
RS_MD5_Uvcc_N        MD4_Inv5_1 com 1G
.MODEL        _MD5_Uvcc_N VSWITCH Roff=1e6 Ron=1 Voff=0.01 Von=4.99
S_MD5_Nand_P1         MD5_Nand_5 MD5_OLS_1 MD4_Inv5_1 VSS _MD5_Nand_P1
RS_MD5_Nand_P1        MD4_Inv5_1 VSS 1G
.MODEL        _MD5_Nand_P1 VSWITCH Roff=1e6 Ron=1 Voff=4.9 Von=0.1
S_MD5_Nand_N1         MD5_OLS_1 MD5_Nand_4 MD3_DlyLS_8 VSS _MD5_Nand_N1
RS_MD5_Nand_N1        MD3_DlyLS_8 VSS 1G
.MODEL        _MD5_Nand_N1 VSWITCH Roff=1e6 Ron=1 Voff=0.1 Von=4.9
S_MD5_Nand_P2         MD5_Nand_5 MD5_OLS_1 MD3_DlyLS_8 VSS _MD5_Nand_P2
RS_MD5_Nand_P2        MD3_DlyLS_8 VSS 1G
.MODEL        _MD5_Nand_P2 VSWITCH Roff=1e6 Ron=1 Voff=4.9 Von=0.1
V_MD5_Nand_V         MD5_Nand_5 VSS 5V
S_MD5_Nand_N2         MD5_Nand_4 VSS MD4_Inv5_1 VSS _MD5_Nand_N2
RS_MD5_Nand_N2        MD4_Inv5_1 VSS 1G
.MODEL        _MD5_Nand_N2 VSWITCH Roff=1e6 Ron=1 Voff=0.1 Von=4.9
S_MD5_OLS_P         VCC MD5_OLS_2 MD5_OLS_1 com _MD5_OLS_P
RS_MD5_OLS_P        MD5_OLS_1 com 1G
.MODEL        _MD5_OLS_P VSWITCH Roff=1e9 Ron=1m Voff=4.9 Von=0.1
S_MD5_OLS_N         MD5_OLS_3 com MD5_OLS_1 com _MD5_OLS_N
RS_MD5_OLS_N        MD5_OLS_1 com 1G
.MODEL        _MD5_OLS_N VSWITCH Roff=1e9 Ron=1m Voff=0.1 Von=4.9
R_MD5_OLS_R6         LO MD5_OLS_2 11.4 TC=0.00190676, 9.3240e-07
R_MD5_OLS_R7         MD5_OLS_3 LO 7.76 TC=0.00241396, 2.331e-06
R_MD5_R         com VCC 83.3k TC=-0.00358599, 0.0000124556
D_MD5_D3         com VCC diode25 
D_MD4_D2         HO VB diode25 
D_MD4_D1         VS VB diode25 
D_MD4_D4         com VB diode625 
D_MD4_D5         com VS diode625 
D_MD4_D3         VS HO diode25 
C_MD4_C3         VS HO  10p IC=0 
C_MD4_Uvbs_c1         MD4_Uvbs_2 MD4_Uvbs_4  10n  
C_MD4_Uvbs_c2         MD4_Uvbs_5 MD4_Uvbs_2  10n  
C_MD4_Uvbs_c3         com MD4_Inv4_1  10p  
E_MD4_Uvbs_ABM18         MD4_Uvbs_4 com   VALUE {
+  V(VS)+8.4+(8.9-8.4)/(125+40)*(TEMP+40)     }
E_MD4_Uvbs_ABM19         MD4_Uvbs_5 com   VALUE {
+  V(VS)+8.0+(8.45-8.0)/(125+40)*(TEMP+40)    }
X_MD4_Uvbs_Comp         VB MD4_Uvbs_2 MD4_Inv4_1 com COMP
S_MD4_Uvbs_P         MD4_Uvbs_4 MD4_Uvbs_2 MD4_Inv4_1 com _MD4_Uvbs_P
RS_MD4_Uvbs_P        MD4_Inv4_1 com 1G
.MODEL        _MD4_Uvbs_P VSWITCH Roff=1e6 Ron=1 Voff=4.99 Von=0.01
S_MD4_Uvbs_N         MD4_Uvbs_2 MD4_Uvbs_5 MD4_Inv4_1 com _MD4_Uvbs_N
RS_MD4_Uvbs_N        MD4_Inv4_1 com 1G
.MODEL        _MD4_Uvbs_N VSWITCH Roff=1e6 Ron=1 Voff=0.01 Von=4.99
V_MD4_Inv3_V         MD4_Inv3_2 VSS 5V
C_MD4_Inv3_C         VSS MD4_OHS_1  1p  
S_MD4_Inv3_P         MD4_Inv3_2 MD4_OHS_1 MD4_RS_4 VSS _MD4_Inv3_P
RS_MD4_Inv3_P        MD4_RS_4 VSS 1G
.MODEL        _MD4_Inv3_P VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD4_Inv3_N         MD4_OHS_1 VSS MD4_RS_4 VSS _MD4_Inv3_N
RS_MD4_Inv3_N        MD4_RS_4 VSS 1G
.MODEL        _MD4_Inv3_N VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
C_MD4_RS_C7         MD4_RS_6 MD4_RS_5  10p  
C_MD4_RS_C2         VSS MD4_Inv2_3  10p IC=0 
C_MD4_RS_C3         VSS MD3_DlyHS_8  10p IC=0 
C_MD4_RS_C10         MD4_RS_7 MD4_RS_5  10p  
C_MD4_RS_C11         MD4_RS_3 MD4_RS_7  10p  
C_MD4_RS_C12         VSS MD4_RS_3  10p  
C_MD4_RS_C9         VSS MD4_RS_4  10p  
C_MD4_RS_C8         MD4_RS_4 MD4_RS_6  10p  
C_MD4_RS_C1         VSS MD4_RS_4  10p IC=0 
S_MD4_RS_P1         MD4_RS_5 MD4_RS_6 MD4_Inv2_3 VSS _MD4_RS_P1
RS_MD4_RS_P1        MD4_Inv2_3 VSS 1G
.MODEL        _MD4_RS_P1 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD4_RS_P2         MD4_RS_6 MD4_RS_4 MD4_RS_3 VSS _MD4_RS_P2
RS_MD4_RS_P2        MD4_RS_3 VSS 1G
.MODEL        _MD4_RS_P2 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD4_RS_N1         MD4_RS_4 VSS MD4_RS_3 VSS _MD4_RS_N1
RS_MD4_RS_N1        MD4_RS_3 VSS 1G
.MODEL        _MD4_RS_N1 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
S_MD4_RS_P3         MD4_RS_5 MD4_RS_7 MD3_DlyHS_8 VSS _MD4_RS_P3
RS_MD4_RS_P3        MD3_DlyHS_8 VSS 1G
.MODEL        _MD4_RS_P3 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD4_RS_P4         MD4_RS_7 MD4_RS_3 MD4_RS_4 VSS _MD4_RS_P4
RS_MD4_RS_P4        MD4_RS_4 VSS 1G
.MODEL        _MD4_RS_P4 VSWITCH Roff=1e6 Ron=1m Voff=4.9V Von=0.1V
S_MD4_RS_N3         MD4_RS_3 VSS MD3_DlyHS_8 VSS _MD4_RS_N3
RS_MD4_RS_N3        MD3_DlyHS_8 VSS 1G
.MODEL        _MD4_RS_N3 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
V_MD4_RS_V1         MD4_RS_5 VSS 5V
S_MD4_RS_N4         MD4_RS_3 VSS MD4_RS_4 VSS _MD4_RS_N4
RS_MD4_RS_N4        MD4_RS_4 VSS 1G
.MODEL        _MD4_RS_N4 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
S_MD4_RS_N2         MD4_RS_4 VSS MD4_Inv2_3 VSS _MD4_RS_N2
RS_MD4_RS_N2        MD4_Inv2_3 VSS 1G
.MODEL        _MD4_RS_N2 VSWITCH Roff=1e8 Ron=1m Voff=0.1V Von=4.9V
V_MD4_Inv2_V         MD4_Inv2_2 VSS 5V
C_MD4_Inv2_C         VSS MD4_Inv2_3  1p  
S_MD4_Inv2_P         MD4_Inv2_2 MD4_Inv2_3 MD4_Nor1_5 VSS _MD4_Inv2_P
RS_MD4_Inv2_P        MD4_Nor1_5 VSS 1G
.MODEL        _MD4_Inv2_P VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD4_Inv2_N         MD4_Inv2_3 VSS MD4_Nor1_5 VSS _MD4_Inv2_N
RS_MD4_Inv2_N        MD4_Nor1_5 VSS 1G
.MODEL        _MD4_Inv2_N VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
V_MD4_Inv1_V         MD4_Inv1_2 VSS 5V
C_MD4_Inv1_C         VSS MD4_Nor1_1  1p  
S_MD4_Inv1_P         MD4_Inv1_2 MD4_Nor1_1 MD3_DlyHS_8 VSS _MD4_Inv1_P
RS_MD4_Inv1_P        MD3_DlyHS_8 VSS 1G
.MODEL        _MD4_Inv1_P VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD4_Inv1_N         MD4_Nor1_1 VSS MD3_DlyHS_8 VSS _MD4_Inv1_N
RS_MD4_Inv1_N        MD3_DlyHS_8 VSS 1G
.MODEL        _MD4_Inv1_N VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
V_MD4_Inv4_V         MD4_Inv4_2 VSS 5V
C_MD4_Inv4_C         VSS MD4_Nor2_2  1p  
S_MD4_Inv4_P         MD4_Inv4_2 MD4_Nor2_2 MD4_Inv4_1 VSS _MD4_Inv4_P
RS_MD4_Inv4_P        MD4_Inv4_1 VSS 1G
.MODEL        _MD4_Inv4_P VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD4_Inv4_N         MD4_Nor2_2 VSS MD4_Inv4_1 VSS _MD4_Inv4_N
RS_MD4_Inv4_N        MD4_Inv4_1 VSS 1G
.MODEL        _MD4_Inv4_N VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
V_MD4_Nor1_V         MD4_Nor1_3 VSS 5V
S_MD4_Nor1_P1         MD4_Nor1_3 MD4_Nor1_4 MD4_Nor1_1 VSS _MD4_Nor1_P1
RS_MD4_Nor1_P1        MD4_Nor1_1 VSS 1G
.MODEL        _MD4_Nor1_P1 VSWITCH Roff=1e6 Ron=1 Voff=4.9 Von=0.1
S_MD4_Nor1_P2         MD4_Nor1_4 MD4_Nor1_5 MD4_Inv6_3 VSS _MD4_Nor1_P2
RS_MD4_Nor1_P2        MD4_Inv6_3 VSS 1G
.MODEL        _MD4_Nor1_P2 VSWITCH Roff=1e6 Ron=1 Voff=4.9 Von=0.1
S_MD4_Nor1_N1         MD4_Nor1_5 VSS MD4_Inv6_3 VSS _MD4_Nor1_N1
RS_MD4_Nor1_N1        MD4_Inv6_3 VSS 1G
.MODEL        _MD4_Nor1_N1 VSWITCH Roff=1e6 Ron=1 Voff=0.1 Von=4.9
S_MD4_Nor1_N2         MD4_Nor1_5 VSS MD4_Nor1_1 VSS _MD4_Nor1_N2
RS_MD4_Nor1_N2        MD4_Nor1_1 VSS 1G
.MODEL        _MD4_Nor1_N2 VSWITCH Roff=1e6 Ron=1 Voff=0.1 Von=4.9
V_MD4_Inv5_V         MD4_Inv5_2 VSS 5V
C_MD4_Inv5_C         VSS MD4_Nor2_1  1p  
S_MD4_Inv5_P         MD4_Inv5_2 MD4_Nor2_1 MD4_Inv5_1 VSS _MD4_Inv5_P
RS_MD4_Inv5_P        MD4_Inv5_1 VSS 1G
.MODEL        _MD4_Inv5_P VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD4_Inv5_N         MD4_Nor2_1 VSS MD4_Inv5_1 VSS _MD4_Inv5_N
RS_MD4_Inv5_N        MD4_Inv5_1 VSS 1G
.MODEL        _MD4_Inv5_N VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
V_MD4_Nor2_V         MD4_Nor2_3 VSS 5V
S_MD4_Nor2_P1         MD4_Nor2_3 MD4_Nor2_4 MD4_Nor2_1 VSS _MD4_Nor2_P1
RS_MD4_Nor2_P1        MD4_Nor2_1 VSS 1G
.MODEL        _MD4_Nor2_P1 VSWITCH Roff=1e6 Ron=1 Voff=4.9 Von=0.1
S_MD4_Nor2_P2         MD4_Nor2_4 MD4_Inv6_1 MD4_Nor2_2 VSS _MD4_Nor2_P2
RS_MD4_Nor2_P2        MD4_Nor2_2 VSS 1G
.MODEL        _MD4_Nor2_P2 VSWITCH Roff=1e6 Ron=1 Voff=4.9 Von=0.1
S_MD4_Nor2_N1         MD4_Inv6_1 VSS MD4_Nor2_2 VSS _MD4_Nor2_N1
RS_MD4_Nor2_N1        MD4_Nor2_2 VSS 1G
.MODEL        _MD4_Nor2_N1 VSWITCH Roff=1e6 Ron=1 Voff=0.1 Von=4.9
S_MD4_Nor2_N2         MD4_Inv6_1 VSS MD4_Nor2_1 VSS _MD4_Nor2_N2
RS_MD4_Nor2_N2        MD4_Nor2_1 VSS 1G
.MODEL        _MD4_Nor2_N2 VSWITCH Roff=1e6 Ron=1 Voff=0.1 Von=4.9
V_MD4_Inv6_V         MD4_Inv6_2 VSS 5V
C_MD4_Inv6_C         VSS MD4_Inv6_3  1p  
S_MD4_Inv6_P         MD4_Inv6_2 MD4_Inv6_3 MD4_Inv6_1 VSS _MD4_Inv6_P
RS_MD4_Inv6_P        MD4_Inv6_1 VSS 1G
.MODEL        _MD4_Inv6_P VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD4_Inv6_N         MD4_Inv6_3 VSS MD4_Inv6_1 VSS _MD4_Inv6_N
RS_MD4_Inv6_N        MD4_Inv6_1 VSS 1G
.MODEL        _MD4_Inv6_N VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
R_MD4_R1         VS VB 120k TC=-0.00135415, -2.516e-7
S_MD4_OHS_P         VB MD4_OHS_2 MD4_OHS_1 com _MD4_OHS_P
RS_MD4_OHS_P        MD4_OHS_1 com 1G
.MODEL        _MD4_OHS_P VSWITCH Roff=1e9 Ron=1m Voff=4.9 Von=0.1
S_MD4_OHS_N         MD4_OHS_3 VS MD4_OHS_1 com _MD4_OHS_N
RS_MD4_OHS_N        MD4_OHS_1 com 1G
.MODEL        _MD4_OHS_N VSWITCH Roff=1e9 Ron=1m Voff=0.1 Von=4.9
R_MD4_OHS_R6         HO MD4_OHS_2 11.4 TC=0.00190676, 9.3240e-07
R_MD4_OHS_R7         MD4_OHS_3 HO 7.76 TC=0.00241396, 2.331e-06
C_MD3_C1         com MD3_DlyHS_8  10p  
C_MD3_C2         com MD3_DlyLS_8  10p  
E_MD3_ABM21         MD3_DlyHS_1 com   VALUE { ( V(VB)  
+ -V(VS) )   }
C_MD3_DlyHS_C         VSS MD3_DlyHS_5  10n  
S_MD3_DlyHS_delay_P         MD3_DlyHS_20 MD3_DlyHS_5 MD3_DlyHS_2 VSS
+  _MD3_DlyHS_delay_P
RS_MD3_DlyHS_delay_P        MD3_DlyHS_2 VSS 1G
.MODEL        _MD3_DlyHS_delay_P VSWITCH Roff=1e6 Ron=10 Voff=4.99V Von=0.01V
S_MD3_DlyHS_delay_N         MD3_DlyHS_5 VSS MD3_DlyHS_2 VSS _MD3_DlyHS_delay_N
RS_MD3_DlyHS_delay_N        MD3_DlyHS_2 VSS 1G
.MODEL        _MD3_DlyHS_delay_N VSWITCH Roff=1e6 Ron=10 Voff=0.01V Von=4.99V
S_MD3_DlyHS_P1         MD3_DlyHS_10 MD3_DlyHS_11 MD3_DlyHS_6 VSS _MD3_DlyHS_P1
RS_MD3_DlyHS_P1        MD3_DlyHS_6 VSS 1G
.MODEL        _MD3_DlyHS_P1 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD3_DlyHS_P2         MD3_DlyHS_11 MD3_DlyHS_9 MD3_DlyHS_8 VSS _MD3_DlyHS_P2
RS_MD3_DlyHS_P2        MD3_DlyHS_8 VSS 1G
.MODEL        _MD3_DlyHS_P2 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD3_DlyHS_N1         MD3_DlyHS_9 VSS MD3_DlyHS_8 VSS _MD3_DlyHS_N1
RS_MD3_DlyHS_N1        MD3_DlyHS_8 VSS 1G
.MODEL        _MD3_DlyHS_N1 VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
S_MD3_DlyHS_MP1         MD3_DlyHS_12 MD3_DlyHS_13 MD3_DlyHS_9 VSS
+  _MD3_DlyHS_MP1
RS_MD3_DlyHS_MP1        MD3_DlyHS_9 VSS 1G
.MODEL        _MD3_DlyHS_MP1 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD3_DlyHS_MP2         MD3_DlyHS_13 MD3_DlyHS_8 MD3_DlyHS_7 VSS _MD3_DlyHS_MP2
RS_MD3_DlyHS_MP2        MD3_DlyHS_7 VSS 1G
.MODEL        _MD3_DlyHS_MP2 VSWITCH Roff=1e6 Ron=1 Voff=4.9 Von=0.1
S_MD3_DlyHS_MN1         MD3_DlyHS_8 VSS MD3_DlyHS_7 VSS _MD3_DlyHS_MN1
RS_MD3_DlyHS_MN1        MD3_DlyHS_7 VSS 1G
.MODEL        _MD3_DlyHS_MN1 VSWITCH Roff=1e6 Ron=1 Voff=0.1 Von=4.9
S_MD3_DlyHS_MN2         MD3_DlyHS_8 VSS MD3_DlyHS_9 VSS _MD3_DlyHS_MN2
RS_MD3_DlyHS_MN2        MD3_DlyHS_9 VSS 1G
.MODEL        _MD3_DlyHS_MN2 VSWITCH Roff=1e6 Ron=1 Voff=0.1 Von=4.9
X_MD3_DlyHS_Comp1         MD3_DlyHS_5 MD3_DlyHS_18 MD3_DlyHS_7 com COMP
X_MD3_DlyHS_Comp2         MD3_DlyHS_3 MD3_DlyHS_5 MD3_DlyHS_6 com COMP
E_MD3_DlyHS_ABM5         MD3_DlyHS_21 com   VALUE { (5-5*EXP(-{toffT2}/10/10n))  
+ *(5-5* EXP(-( {toffT1}+({toffT3}-{toffT1})/({T3}-{T1})*(TEMP-{T1}))/10/10n))
+   
+ /(5-5* EXP(-( {toffT1}+({toffT3}-{toffT1})/({T3}-{T1})*({T2}-{T1}))/10/10n))
+   }
E_MD3_DlyHS_ABM14         MD3_DlyHS_19 com   VALUE { (1-EXP(-( {toffVdd1}+(
+ {toffVdd3}-{toffVdd1})/({V3}-{V1})*(V(VDD)-{V1}))/10/ 10n))/  
+ (1-EXP(-( {toffVdd1}+({toffVdd3}-{toffVdd1})/({V3}-{V1})*({V2}  -{V1}))/10/
+  10n))   }
E_MD3_DlyHS_ABM31         MD3_DlyHS_18 com   VALUE { ( V(MD3_DlyHS_21)  
+ *V(MD3_DlyHS_17)  
+ *V(MD3_DlyHS_19) )   }
E_MD3_DlyHS_ABM24         MD3_DlyHS_3 com   VALUE { (EXP(-({tonVdd1}+({tonVdd3}-
+ {tonVdd1})/({V3}-{V1})*(V(VDD)-{V1}))/10/10n))/((EXP(-({tonVdd1}+({tonVdd3}-
+ {tonVdd1})/({V3}-{V1})*({V2}-  {V1}))/10/10n)))  
+ *(5* EXP(-( {tonT1}+({tonT3}-{tonT1})/({T3}-{T1})*(TEMP-{T1})) /10/
+  10n))/(5* EXP(-( {tonT1}+({tonT3}-{tonT1})/({T3}-{T1})*({T2}-{T1})) /10/
+  10n))*5*EXP(-{tonT2}/10/10n)* (EXP(-({tonV1}+({tonV3}-{tonV1})/({V3}-
+ {V1})*(V(MD3_DlyHS_1)-{V1}))/10/10n))/((EXP(-( {tonV1}+({tonV3}-{tonV1})/({V3}-
+ {V1})*({V2}-{V1}))/10/10n)))   }
V_MD3_DlyHS_V_delay         MD3_DlyHS_20 VSS 5V
C_MD3_DlyHS_C3         VSS MD3_DlyHS_6  10p  
V_MD3_DlyHS_VCC1         MD3_DlyHS_10 VSS 5V
C_MD3_DlyHS_C6         VSS MD3_DlyHS_9  10p IC=-5V 
C_MD3_DlyHS_C5         VSS MD3_DlyHS_8  10p IC=0V 
V_MD3_DlyHS_VCC2         MD3_DlyHS_12 VSS 5V
S_MD3_DlyHS_N2         MD3_DlyHS_9 VSS MD3_DlyHS_6 VSS _MD3_DlyHS_N2
RS_MD3_DlyHS_N2        MD3_DlyHS_6 VSS 1G
.MODEL        _MD3_DlyHS_N2 VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
C_MD3_DlyHS_C4         VSS MD3_DlyHS_7  10p  
E_MD3_DlyHS_ABM13         MD3_DlyHS_17 com   VALUE { (1-EXP(-( {toffV1}+({toffV3}-
+ {toffV1})/({V3}-{V1})*((V(MD3_DlyHS_1))-{V1}))/10/ 10n))/  
+ (1-EXP(-( {toffV1}+({toffV3}-{toffV1})/({V3}-{V1})*({V2}  -{V1}))/10/ 10n)) 
+   }
C_MD3_DlyLS_C         VSS MD3_DlyLS_5  10n  
S_MD3_DlyLS_delay_P         MD3_DlyLS_20 MD3_DlyLS_5 MD3_DlyLS_2 VSS
+  _MD3_DlyLS_delay_P
RS_MD3_DlyLS_delay_P        MD3_DlyLS_2 VSS 1G
.MODEL        _MD3_DlyLS_delay_P VSWITCH Roff=1e6 Ron=10 Voff=4.99V Von=0.01V
S_MD3_DlyLS_delay_N         MD3_DlyLS_5 VSS MD3_DlyLS_2 VSS _MD3_DlyLS_delay_N
RS_MD3_DlyLS_delay_N        MD3_DlyLS_2 VSS 1G
.MODEL        _MD3_DlyLS_delay_N VSWITCH Roff=1e6 Ron=10 Voff=0.01V Von=4.99V
S_MD3_DlyLS_P1         MD3_DlyLS_10 MD3_DlyLS_11 MD3_DlyLS_6 VSS _MD3_DlyLS_P1
RS_MD3_DlyLS_P1        MD3_DlyLS_6 VSS 1G
.MODEL        _MD3_DlyLS_P1 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD3_DlyLS_P2         MD3_DlyLS_11 MD3_DlyLS_9 MD3_DlyLS_8 VSS _MD3_DlyLS_P2
RS_MD3_DlyLS_P2        MD3_DlyLS_8 VSS 1G
.MODEL        _MD3_DlyLS_P2 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD3_DlyLS_N1         MD3_DlyLS_9 VSS MD3_DlyLS_8 VSS _MD3_DlyLS_N1
RS_MD3_DlyLS_N1        MD3_DlyLS_8 VSS 1G
.MODEL        _MD3_DlyLS_N1 VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
S_MD3_DlyLS_MP1         MD3_DlyLS_12 MD3_DlyLS_13 MD3_DlyLS_9 VSS
+  _MD3_DlyLS_MP1
RS_MD3_DlyLS_MP1        MD3_DlyLS_9 VSS 1G
.MODEL        _MD3_DlyLS_MP1 VSWITCH Roff=1e6 Ron=1 Voff=4.9V Von=0.1V
S_MD3_DlyLS_MP2         MD3_DlyLS_13 MD3_DlyLS_8 MD3_DlyLS_7 VSS _MD3_DlyLS_MP2
RS_MD3_DlyLS_MP2        MD3_DlyLS_7 VSS 1G
.MODEL        _MD3_DlyLS_MP2 VSWITCH Roff=1e6 Ron=1 Voff=4.9 Von=0.1
S_MD3_DlyLS_MN1         MD3_DlyLS_8 VSS MD3_DlyLS_7 VSS _MD3_DlyLS_MN1
RS_MD3_DlyLS_MN1        MD3_DlyLS_7 VSS 1G
.MODEL        _MD3_DlyLS_MN1 VSWITCH Roff=1e6 Ron=1 Voff=0.1 Von=4.9
S_MD3_DlyLS_MN2         MD3_DlyLS_8 VSS MD3_DlyLS_9 VSS _MD3_DlyLS_MN2
RS_MD3_DlyLS_MN2        MD3_DlyLS_9 VSS 1G
.MODEL        _MD3_DlyLS_MN2 VSWITCH Roff=1e6 Ron=1 Voff=0.1 Von=4.9
X_MD3_DlyLS_Comp1         MD3_DlyLS_5 MD3_DlyLS_18 MD3_DlyLS_7 com COMP
X_MD3_DlyLS_Comp2         MD3_DlyLS_3 MD3_DlyLS_5 MD3_DlyLS_6 com COMP
E_MD3_DlyLS_ABM5         MD3_DlyLS_21 com   VALUE { (5-5*EXP(-{toffT2}/10/10n))  
+ *(5-5* EXP(-( {toffT1}+({toffT3}-{toffT1})/({T3}-{T1})*(TEMP-{T1}))/10/10n))
+   
+ /(5-5* EXP(-( {toffT1}+({toffT3}-{toffT1})/({T3}-{T1})*({T2}-{T1}))/10/10n))
+   }
E_MD3_DlyLS_ABM14         MD3_DlyLS_19 com   VALUE { (1-EXP(-( {toffVdd1}+(
+ {toffVdd3}-{toffVdd1})/({V3}-{V1})*(V(VDD)-{V1}))/10/ 10n))/  
+ (1-EXP(-( {toffVdd1}+({toffVdd3}-{toffVdd1})/({V3}-{V1})*({V2}  -{V1}))/10/
+  10n))   }
E_MD3_DlyLS_ABM31         MD3_DlyLS_18 com   VALUE { ( V(MD3_DlyLS_21)  
+ *V(MD3_DlyLS_17)  
+ *V(MD3_DlyLS_19) )   }
E_MD3_DlyLS_ABM24         MD3_DlyLS_3 com   VALUE { (EXP(-({tonVdd1}+({tonVdd3}-
+ {tonVdd1})/({V3}-{V1})*(V(VDD)-{V1}))/10/10n))/((EXP(-({tonVdd1}+({tonVdd3}-
+ {tonVdd1})/({V3}-{V1})*({V2}-  {V1}))/10/10n)))  
+ *(5* EXP(-( {tonT1}+({tonT3}-{tonT1})/({T3}-{T1})*(TEMP-{T1})) /10/
+  10n))/(5* EXP(-( {tonT1}+({tonT3}-{tonT1})/({T3}-{T1})*({T2}-{T1})) /10/
+  10n))*5*EXP(-{tonT2}/10/10n)* (EXP(-({tonV1}+({tonV3}-{tonV1})/({V3}-
+ {V1})*(V(VCC)-{V1}))/10/10n))/((EXP(-( {tonV1}+({tonV3}-{tonV1})/({V3}-{V1})*(
+ {V2}-{V1}))/10/10n)))   }
V_MD3_DlyLS_V_delay         MD3_DlyLS_20 VSS 5V
C_MD3_DlyLS_C3         VSS MD3_DlyLS_6  10p  
V_MD3_DlyLS_VCC1         MD3_DlyLS_10 VSS 5V
C_MD3_DlyLS_C6         VSS MD3_DlyLS_9  10p IC=-5V 
C_MD3_DlyLS_C5         VSS MD3_DlyLS_8  10p IC=0V 
V_MD3_DlyLS_VCC2         MD3_DlyLS_12 VSS 5V
S_MD3_DlyLS_N2         MD3_DlyLS_9 VSS MD3_DlyLS_6 VSS _MD3_DlyLS_N2
RS_MD3_DlyLS_N2        MD3_DlyLS_6 VSS 1G
.MODEL        _MD3_DlyLS_N2 VSWITCH Roff=1e6 Ron=1 Voff=0.1V Von=4.9V
C_MD3_DlyLS_C4         VSS MD3_DlyLS_7  10p  
E_MD3_DlyLS_ABM13         MD3_DlyLS_17 com   VALUE { (1-EXP(-( {toffV1}+({toffV3}-
+ {toffV1})/({V3}-{V1})*((V(VCC))-{V1}))/10/ 10n))/  
+ (1-EXP(-( {toffV1}+({toffV3}-{toffV1})/({V3}-{V1})*({V2}  -{V1}))/10/ 10n)) 
+   }

.ENDS    IR2113

.SUBCKT COMP 1 2 3 4
E1 5 4 VALUE={IF((V(1)>V(2)), V(4)+5V, V(4))}
R1 5 3 1
C1 3 4 10P
.ENDS

* SPICE netlist written by S-Edit Win32 11.40
* Written on Sep 5, 2013 at 12:29:29

.SUBCKT BUFFER_2736_5040 IN OUTN OUTP Vminus Vplus
MN1 N25 IN Vminus Vminus NCH W=60u L=4u M=4 AS=0p PS=0u AD=198p PD=52u
MN2 N27 N25 Vminus Vminus NCH W=68u L=4u M=12 AS=0p PS=0u AD=254p PD=60u
MN3 OUTN N27 Vminus Vminus NCH W=76u L=4u M=36 AS=0p PS=0u AD=310p PD=68u
MP1 N26 IN Vplus Vplus PCH W=54u L=4u M=8 AS=0p PS=0u AD=150p PD=45u
MP2 N28 N26 Vplus Vplus PCH W=62u L=4u M=24 AS=0p PS=0u AD=198p PD=53u
MP3 OUTP N28 Vplus Vplus PCH W=70u L=4u M=72 AS=0p PS=0u AD=246p PD=61u
R1 N25 N26  RES 11.7k
R2 N27 N28  RES 1k
R3 OUTN OUTP  RES 100
.ENDS

.SUBCKT espdIN2 A Y COM Vcc
D1 A Vcc DIODE AREA=1378e-12 M=1
D2 COM A DIODE AREA=1322e-12 M=1
D3 COM Y DIODE AREA=630e-12 M=1
MN1 Y COM COM COM NCH W=154u L=4u M=2 AS=0p PS=0u AD=836p PD=143u
R1 Y A  RES 96
.ENDS

.SUBCKT espdIN A Y COM
D1 COM A DIODE AREA=1296e-12 M=1
D2 COM Y DIODE AREA=630e-12 M=1
MN1 Y COM COM COM NCH W=154u L=4u M=2 AS=0p PS=0u AD=836p PD=143u
R1 Y A  RES 96
.ENDS

.SUBCKT espdOUT A COM Vcc
D1 A Vcc DIODE AREA=2806e-12 M=1
D2 COM A DIODE AREA=2000e-12 M=1
.ENDS

.SUBCKT espdOUT_VSVB A VB VS
D1 A VB DIODE AREA=2806e-12 M=1
D2 VS A DIODE AREA=1490e-12 M=1
.ENDS

.SUBCKT INV_60_108 A Y COM Vcc
MN1 Y A COM COM NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MP1 Y A Vcc Vcc PCH W=54u L=4u M=2 AS=0p PS=0u AD=150p PD=45u
.ENDS

.SUBCKT INV_60_108_VSVB A VB VS Y
MN1 Y A VS VS NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MP1 Y A VB VB PCH W=54u L=4u M=2 AS=0p PS=0u AD=150p PD=45u
.ENDS

.SUBCKT LRS NRES NSET QN Vminus Vplus
MN1 p2 p3 N5 Vminus NCH W=60u L=4u M=1 AS=1490p PS=256u AD=198p PD=52u
MN2 N5 NSET Vminus Vminus NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN3 N9 p1 N13 Vminus NCH W=60u L=4u M=1 AS=1490p PS=256u AD=198p PD=52u
MN4 N13 NRES Vminus Vminus NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN5 N9 p1 N21 Vminus NCH W=60u L=4u M=1 AS=1490p PS=256u AD=198p PD=52u
MN6 N21 NRES Vminus Vminus NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN7 QN p2 Vminus Vminus NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MP1 p1 NSET Vplus Vplus PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP2 p1 p3 Vplus Vplus PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP3 p3 NRES Vplus Vplus PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP4 p3 p1 Vplus Vplus PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP5 QN p1 Vplus Vplus PCH W=54u L=4u M=2 AS=0p PS=0u AD=150p PD=45u
R1 p2 p1  RES 5k
R2 N9 p3  RES 5k
.ENDS

.SUBCKT NAND2_30_54 A B Y COM Vcc
MN1 Y A N3 COM NCH W=60u L=4u M=1 AS=1490p PS=256u AD=198p PD=52u
MN2 N3 B COM COM NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN3 Y B N10 COM NCH W=60u L=4u M=1 AS=1490p PS=256u AD=198p PD=52u
MN4 N10 A COM COM NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MP1 Y A Vcc Vcc PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP2 Y B Vcc Vcc PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
.ENDS

.SUBCKT NOR2_60_54 A B Y COM Vcc
MN1 Y A COM COM NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN2 Y B COM COM NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MP1 N11 A Vcc Vcc PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP2 Y B N11 Vcc PCH W=54u L=4u M=1 AS=1058p PS=183u AD=150p PD=45u
MP3 N18 B Vcc Vcc PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP4 Y A N18 Vcc PCH W=54u L=4u M=1 AS=1058p PS=183u AD=150p PD=45u
.ENDS

.SUBCKT NOR2_60_54_VSVB A B VB VS Y
MN1 Y A VS VS NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN2 Y B VS VS NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MP1 N11 A VB VB PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP2 Y B N11 VB PCH W=54u L=4u M=1 AS=1058p PS=183u AD=150p PD=45u
MP3 N18 B VB VB PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP4 Y A N18 VB PCH W=54u L=4u M=1 AS=1058p PS=183u AD=150p PD=45u
.ENDS

.SUBCKT TSH A Y COM Vcc
MN1 Y A N3 COM NCH W=60u L=4u M=1 AS=1490p PS=256u AD=198p PD=52u
MN2 N3 A COM COM NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN3 Vcc Y N3 COM NCH W=60u L=4u M=1 AS=1490p PS=256u AD=198p PD=52u
MP1 N15 A Vcc Vcc PCH W=54u L=4u M=2 AS=0p PS=0u AD=150p PD=45u
MP2 Y A N15 Vcc PCH W=54u L=4u M=2 AS=1058p PS=183u AD=150p PD=45u
MP3 COM Y N15 Vcc PCH W=54u L=4u M=2 AS=1058p PS=183u AD=150p PD=45u
.ENDS

.SUBCKT UV_Detector OUT Vminus Vplus
C1 N1 Vminus CAP 5pF M=2
C2 N20 Vminus CAP 5pF M=1
C3 N20 Vminus CAP 2pF M=1
MN1 N16 N16 Vminus Vminus NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN2 s1 N1 N15 Vminus NCH W=60u L=4u M=2 AS=1490p PS=256u AD=198p PD=52u
MN3 N15 N16 Vminus Vminus NCH W=60u L=4u M=8 AS=0p PS=0u AD=198p PD=52u
MN4 s2 N20 N15 Vminus NCH W=60u L=4u M=2 AS=1490p PS=256u AD=198p PD=52u
MN5 N28 N28 Vminus Vminus NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN6 N76 N28 Vminus Vminus NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN7 OUT N76 Vminus Vminus NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MP1 N16 N16 N1 Vplus PCH W=54u L=4u M=1 AS=1058p PS=183u AD=150p PD=45u
MP2 s1 s1 Vplus Vplus PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP3 s1 s2 Vplus Vplus PCH W=100u L=4u M=1 AS=0p PS=0u AD=426p PD=91u
MP4 s2 s1 Vplus Vplus PCH W=100u L=4u M=1 AS=0p PS=0u AD=426p PD=91u
MP5 s2 s2 Vplus Vplus PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP6 N28 s1 Vplus Vplus PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP7 N61 s2 Vplus Vplus PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP8 OUT N61 Vplus Vplus PCH W=54u L=4u M=2 AS=0p PS=0u AD=150p PD=45u
R1 N1 Vplus  RES 711.7k
R2 N69 Vplus  RES 425k
R3 N71 N69  RES 40k
R4 N20 N71  RES 20k
R5 N73 N20  RES 30k
R6 N74 N73  RES 30k
R7 Vminus N74  RES 315k
R8 N76 N61  RES 6.8k
.ENDS

* Main circuit: TopLevel
XBUFFER_2736_5040_1 N52 N89 N76 VS VB BUFFER_2736_5040
XBUFFER_2736_5040_2 N63 N90 N92 COM Vcc BUFFER_2736_5040
C1 N68 COM CAP 2pF M=4
C2 Vcc COM CAP 5pF M=6
C3 Vcc COM CAP 2pF M=1
C4 Vcc COM CAP 1pF M=13
C5 N74 COM CAP 1pF M=3
C6 N77 N78 CAP 22.8pF M=1
C7 N78 N75 CAP 22.8pF M=1
C8 N75 s1 CAP 22.8pF M=1
C9 N81 N82 CAP 22.8pF M=1
C10 N82 N79 CAP 22.8pF M=1
C11 N79 s2 CAP 22.8pF M=1
D1 COM Vcc DIODE AREA=2215e-12 M=1
D2 COM Vcc DIODE AREA=2806e-12 M=1
D3 s1 Vcc DIODE AREA=1000e-12 M=1
D4 s2 Vcc DIODE AREA=1000e-12 M=1
D5 VS VB DIODE AREA=2806e-12 M=1
D6 VS VB DIODE AREA=1000e-12 M=1
D7 VS VB DIODE AREA=1492e-12 M=1
D8 p1 VB DIODE AREA=2000e-12 M=1
D9 VS p1 DIODE AREA=2000e-12 M=1
D10 p2 VB DIODE AREA=2000e-12 M=1
D11 VS p2 DIODE AREA=2000e-12 M=1
XespdIN2_1 CX N68 COM Vcc espdIN2
XespdIN_1 IN N71 COM espdIN
XespdOUT_1 LO COM Vcc espdOUT
XespdOUT_VSVB_1 HO VB VS espdOUT_VSVB
XINV_60_108_1 N6 N70 COM Vcc INV_60_108
XINV_60_108_2 N11 N65 COM Vcc INV_60_108
XINV_60_108_3 N65 N91 COM Vcc INV_60_108
XINV_60_108_4 N67 N63 COM Vcc INV_60_108
XINV_60_108_VSVB_4 x2 VB VS N57 INV_60_108_VSVB
XINV_60_108_VSVB_5 x1 VB VS N55 INV_60_108_VSVB
XINV_60_108_VSVB_6 N55 VB VS N54 INV_60_108_VSVB
XLRS_2 N54 N53 N52 VS VB LRS
MN1 N87 N87 VS VS NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN2 p4 N87 VS VS NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN3 N83 N83 VS VS NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN4 p3 N83 VS VS NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN5 x1 p3 VS VS NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN6 x2 p4 VS VS NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN7 Vcc COM COM COM NCH W=60u L=4u M=8 AS=0p PS=0u AD=198p PD=52u
MN8 s1 N91 COM COM NCH W=60u L=4u M=2 AS=0p PS=0u AD=198p PD=52u
MN9 s2 N65 COM COM NCH W=60u L=4u M=2 AS=0p PS=0u AD=198p PD=52u
MN10 VB VS VS VS NCH W=60u L=4u M=8 AS=0p PS=0u AD=198p PD=52u
MN11 HO N89 VS VS NCH W=80u L=4u M=128 AS=0p PS=0u AD=338p PD=72u
MN12 LO N90 COM COM NCH W=80u L=4u M=128 AS=0p PS=0u AD=338p PD=72u
MN_12 p1 VS VS VS NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MN_13 p2 VS VS VS NCH W=60u L=4u M=1 AS=0p PS=0u AD=198p PD=52u
MP1 N80 N80 VB VB PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP2 N84 N80 VB VB PCH W=54u L=4u M=2 AS=0p PS=0u AD=150p PD=45u
MP3 N87 N72 N84 VB PCH W=54u L=4u M=4 AS=1058p PS=183u AD=150p PD=45u
MP4 p4 N85 N84 VB PCH W=54u L=4u M=4 AS=1058p PS=183u AD=150p PD=45u
MP5 N83 N85 N84 VB PCH W=54u L=4u M=4 AS=1058p PS=183u AD=150p PD=45u
MP6 p3 N72 N84 VB PCH W=54u L=4u M=4 AS=1058p PS=183u AD=150p PD=45u
MP7 x1 x2 VB VB PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP8 x2 x1 VB VB PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP9 N66 N66 VB VB PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP10 N86 N86 VB VB PCH W=54u L=4u M=1 AS=0p PS=0u AD=150p PD=45u
MP11 p1 p1 N66 VB PCH W=54u L=4u M=1 AS=1058p PS=183u AD=150p PD=45u
MP12 p2 p2 N86 VB PCH W=54u L=4u M=1 AS=1058p PS=183u AD=150p PD=45u
MP13 s1 N91 Vcc Vcc PCH W=54u L=4u M=4 AS=0p PS=0u AD=150p PD=45u
MP14 s2 N65 Vcc Vcc PCH W=54u L=4u M=4 AS=0p PS=0u AD=150p PD=45u
MP15 HO N76 VB VB PCH W=74u L=4u M=256 AS=0p PS=0u AD=270p PD=65u
MP16 LO N92 Vcc Vcc PCH W=74u L=4u M=256 AS=0p PS=0u AD=270p PD=65u
XNAND2_30_54_1 N7 N6 N3 COM Vcc NAND2_30_54
XNOR2_60_54_1 N6 N7 N4 COM Vcc NOR2_60_54
XNOR2_60_54_2 N4 N5 N11 COM Vcc NOR2_60_54
XNOR2_60_54_3 N5 N3 N69 COM Vcc NOR2_60_54
XNOR2_60_54_VSVB_2 N56 N57 VB VS N53 NOR2_60_54_VSVB
R1 VS N80  RES 240k
R2 COM N71  RES 500k
R3 N68 N70  RES 67k
R4 N85 p1  RES 1k
R5 N72 p2  RES 1k
R6 N74 N69  RES 15k
R7 N77 p1  RES 5k
R8 N78 N77  RES 333k
R9 N75 N78  RES 333k
R10 s1 N75  RES 333k
R11 N81 p2  RES 5k
R12 N82 N81  RES 333k
R13 N79 N82  RES 333k
R14 s2 N79  RES 333k
XTSH_1 N71 N6 COM Vcc TSH
XTSH_2 N68 N7 COM Vcc TSH
XTSH_3 N74 N67 COM Vcc TSH
XUV_Detector_1 N5 COM AVDD UV_Detector
XUV_Detector_3 N56 VS VB UV_Detector
* End of main circuit: TopLevel

*may2004
*Models for 3u Exiton RING CMOS TRS  
.MODEL NCH NMOS LEVEL=3
+ VTO=0.9
+ UO=400
+ TOX=600e-10
+ LD=0.1e-6
+ WD=0
+ GAMMA=0.045
+ NSUB=1e15
+ PHI=0.7
+ PB=0.9
+ CJ=6e-04
+ CJSW=4.5e-10
+ MJ=0.5
+ MJSW=0.3
+ KF=1
+ AF=1
+ RSH=170
+ XJ=1e-07
+ FC=0.5
+ DELTA=0.1
+ VMAX=1.2e5
+ JS=1.2e-06
+ IS=1e-13
+ ETA=1e-02
+ THETA=2e-2
+ KAPPA=0.3
+ CGSO=4e-10
+ CGDO=4e-10
+ CGBO=22e-10

.MODEL PCH PMOS LEVEL=3
+ VTO=-1.4
+ UO=200
+ TOX=600e-10
+ LD=0.1e-6
+ WD=0
+ GAMMA=0.015
+ NSUB=1e14
+ PHI=0.7
+ PB=0.8
+ CJ=5e-04
+ CJSW=3.5e-10
+ MJ=0.5
+ MJSW=0.3
+ KF=1
+ AF=1
+ RSH=1700
+ XJ=1e-07
+ FC=0.5
+ DELTA=0.1
+ VMAX=1e5
+ JS=1.2e-06
+ IS=1e-13
+ ETA=1e-02
+ THETA=2e-2
+ KAPPA=0.3
+ CGSO=4e-10
+ CGDO=4e-10
+ CGBO=26e-10

.MODEL RES R
+TC1=0.00065

.MODEL CAP C
*+TC1=0.01
*+VC1=0.1

.MODEL DIODE D LEVEL=1
+IS=6e-14
*+RS=10e-12
+N=1.1
+TT=2e-9
+CJO=1e-12
*+CJO=1e-12
+VJ=0.65
*+M=0.4
+FC=0.5
+EG=1.11
+XTI=3
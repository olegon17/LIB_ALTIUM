* TLE2141 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.03 ON 08/15/90 AT 15:59
* REV (N/A)      SUPPLY VOLTAGE: 5V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TLE2141  1 2 3 4 5
*
  C1   11 12 9.741E-12
  C2    6  7 30.00E-12
  C3 87 0 45E-9
  CPSR 85 86 2.65E-9
  DCM+ 81 82 DX
  DCM- 83 81 DX
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  ECMR 84 99 (2,99) 1
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  EPSR 85 0 POLY(1) (3,4) -331E-6 66.2E-6
  ENSE 89 2 POLY(1) (88,0) 225E-6 1
  FB 7 99 POLY(6) VB VC VE VLP VLN VPSR 0 11.62E6 -10E6 10E6 10E6 -10E6 11E6
  GA    6  0 11 12 1.282E-3
  GCM   0  6 10 99 1.614E-9
  GPSR 85 86 (85,86) 100E-6
  GRC1 4 11 (4,11) 1.282E-3
  GRC2 4 12 (4,12) 1.282E-3
  GRE1 13 10 (13,10) 1.349E-3
  GRE2 14 10 (14,10) 1.349E-3
  HLIM 90  0 VLIM 1K
  HCMR 80 1 POLY(2) VCM+ VCM- 0 1E2 1E2
  IRP 3 4 2.048E-3
  IEE   3 10 DC 1.352E-3
  IIO 2 0 8E-9
  I1 88 0 1E-21
  Q1   11  89 13 QX
  Q2   12  80 14 QX
  R2    6  9 100.0E3
  RCM 84 81 1K
  REE  10 99 148.0E3
  RN1 87 0 60E6
  RN2 87 88 6.65E3
  RO1   8  5 15
  RO2   7 99 15
  VCM+ 82 99  .09
  VCM- 83 99 -2.07
  VB    9  0 DC 0
  VC 3 53 DC 1.730
  VE   54  4 DC .8
  VLIM  7  8 DC 0
  VLP  91  0 DC 31
  VLN   0 92 DC 31
  VPSR 0 86 DC 0
.MODEL DX D(IS=800.0E-18)
.MODEL QX PNP(IS=800.0E-18 BF=843.8)
.ENDS

*   SPICE3
.subckt 1N4007 1 2
ddio 1 2 D1n4007

.MODEL D1n4007 d
+IS=7.02767e-09 RS=0.0341512 N=1.80803 EG=1.05743
+XTI=5 BV=1000 IBV=5e-08 CJO=1e-11
+VJ=0.7 M=0.5 FC=0.5 TT=1e-07
+KF=0 AF=1

.ends
* PSpice Model Editor - Version 16.0.0
*****************************************************************************
* (C) Copyright 2009 Texas Instruments Incorporated. All rights reserved.                                            
*****************************************************************************
* Final 2.00
* Changed encrypted model to unencrypted.
*****************************************************************************
.SUBCKT TL431 7 6 11
*             K A FDBK
V1 1 6 2.495
R1 6 2 15.6
C1 2 6 .5U
R2 2 3 100
C2 3 4 .08U
R3 4 6 10
GB1 6 8 VALUE = {IF(V(3,6)< 0 , 1.73*V(3,6) -1U , -1U)}
D1 5 8 DCLAMP
D2 7 8 DCLAMP
V4 5 6 2
G1 6 2 1 11 0.11
.MODEL DCLAMP D (IS=13.5N RS=25M N=1.59
+ CJO=45P VJ=.75 M=.302 TT=50.4N BV=34V IBV=1MA)
.ENDS
*June 23, 2010
*Doc. ID: 90123, Rev. A
*File Name: irfp460n_PS.txt and irfp460n _PS.spi
*This document is intended as a SPICE modeling guideline and does not
*constitute a commercial product data sheet.  Designers should refer to the
*appropriate data sheet of the same number for guaranteed specification
*limits.
.SUBCKT IRFP460 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Aug 23, 01
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=5.44745 LAMBDA=0 KP=6.90602
+CGSO=3.48293e-05 CGDO=1e-12
RS 8 3 0.0001
D1 3 1 MD
.MODEL MD D IS=3.79465e-10 RS=0.0070727 N=1.23149 BV=500
+IBV=0.00025 EG=1.2 XTI=4 TT=0
+CJO=3.99547e-09 VJ=1.87709 M=0.9 FC=0.5
RDS 3 1 1e+06
RD 9 1 0.196416
RG 2 7 2.48359
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=2.45097e-09 VJ=0.904484 M=0.9 FC=1.00001e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=0.403203 RS=3.00029e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 3.43526e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.403203
.ENDS IRFP460

.subckt IR2153 Vcc Rt Ct COM LO VS HO VB 
R5 ARB3_N1 Rt 100 
Rdead ARB3_N2 ARB4_OUT 1k 
Cdead ARB3_N2 COM 1.8n 
RdlyH CdlyH_P ARB5_OUT 1k 
CdlyH CdlyH_P COM 910p 
RdlyL CdlyL_P ARB3_OUT 1k 
CdlyL CdlyL_P COM 910p 
GARB1 Vcc COM VALUE={(75u+500u*(V(Vcc,COM)>8)+5m*exp(10*(V(Vcc,COM)-15.6)))*(V(Vcc,COM)>1)} 
*Micropower startup VCC supply current 75u ; Quiescent VCC supply current 500u; VCC zener clamp voltage 15.6V On ICC = 5mA 
EARB2 ARB3_N1 COM VALUE={V(ARB7_N1,COM)*((V(Ct,COM)<V>4) OR (V(Ct,COM)<V(ARB7_N1,COM)/3 AND V(ARB3_N1,COM)<3>8 AND V(ARB3_N2,COM)>2.5 )* (V(ARB3_N3,COM)>2.5)} 
EARB4 ARB4_OUT COM VALUE={5*( V(ARB3_N1,COM)>0.1 AND V(Ct,COM)>V(ARB3_N1,COM)/3)} 
EARB5 ARB5_OUT COM VALUE={5*( V(ARB3_N1,COM)<8 AND V(ARB3_N2,COM)<2>1)} 
EARB6 ARB7_N1 COM VALUE={V(Vcc,COM)*((V(Vcc,COM)>8 AND V(ARB7_N1,COM)>0.2)OR(V(Vcc,COM)>9 AND V(ARB7_N1,COM)<0>V(ARB7_N1,COM)/6)} ; * for Inhibit LO in SD mode 
GARB8 Ct COM VALUE={(V(ARB7_N1,COM)<1>0.1)} ;* ICTUV UV-mode CT pin pulldown current 0.8mA 
S1 HO VS CdlyH_P COM SVL 
S2 VB HO CdlyH_P COM SVH 
S3 Vcc LO CdlyL_P COM SVH 
S4 LO COM CdlyL_P COM SVL 
.MODEL SVH VSWITCH (RON=50 ROFF=1Meg VON=2.5 VOFF=2.45) 
.MODEL SVL VSWITCH (RON=50 ROFF=1Meg VON=2.45 VOFF=2.5) 
.ends IR2153
*******************************************
*BZV55-C43
*NXP Semiconductors
*
*IR    = 50nA  @ VR   = 0,7V
*IZSM  = 0,6A  @ tp   = 100�s
*VZmax = 46,0V @ IZ   = 2mA
*VZSM  =       @ IZSM =
*
*Package: SOD80C
*
*Package Pin 1: Cathode      
*Package Pin 2: Anode
*
*Simulator: SPICE2
*******************************************
*#
.SUBCKT BZV55C43 1 2
*
*The resistor R1 and the diode D2 do not reflect 
*physical devices but improve 
*only modeling in the reverse 
*mode of operation.
*
R1 1 2 5E+011
D1 1 2 DIODE1
D2 1 2 DIODE2
*
.MODEL DIODE1 D
+ IS = 2E-012
+ N = 1.35
+ BV = 42.17
+ IBV = 6.51E-010
+ RS = 0.5
+ CJO = 1.661E-011
+ VJ = 0.68
+ M = 0.36
+ FC = 0.5
+ TT = 0
+ EG = 1.1
+ XTI = 3
.MODEL DIODE2 D
+ IS = 8.6E-013
+ N = 1.25
+ RS = 5E+005
.ENDS

